/*
*
* Copyright (c) 2013 fpgaminer@bitcoin-mining.com
*
*
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published by
* the Free Software Foundation, either version 3 of the License, or
* (at your option) any later version.
*
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
*
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <http://www.gnu.org/licenses/>.
* 
*/

module vanity_compare (
	input clk,
	input rx_reset,
	input [159:0] rx_min,
	input [159:0] rx_max,
	input [159:0] rx_hash,
	output reg tx_match = 1'b0
);

	always @ (posedge clk)
	begin
		tx_match <= 1'b0;

		if (rx_reset && rx_hash >= rx_min && rx_hash <= rx_max)
			tx_match <= 1'b1;
	end

endmodule
